/****************************************************************************
 * vmon_client_uvm_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: vmon_client_uvm_pkg
 * 
 * TODO: Add package documentation
 */
package vmon_client_uvm_pkg;
	import uvm_pkg::*;
	import vmon_client_pkg::*;

	`include "vmon_client_agent.svh"

endpackage


