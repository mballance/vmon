
/****************************************************************************
 * sv_stub_test_pkg.sv
 ****************************************************************************/

  
/**
 * Package: sv_stub_test_pkg
 * 
 * TODO: Add package documentation
 */
package sv_stub_test_pkg;
	import vmon_bus_monitor_api_pkg::*;
	import vmon_monitor_pkg::*;
	import vmon_client_pkg::*;

	`include "sv_stub_bus_monitor_api.svh"
	`include "sv_stub_test_m2h_path.svh"
	`include "sv_stub_test.svh"


endpackage


